//James Kaden Cassidy jkc.cassidy@gmail.com 12/27/2025

`include "parameters.svh"

module ZIHPM #(

    ) (

    );


endmodule
