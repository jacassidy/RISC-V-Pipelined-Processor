`ifndef GLOBALS_SVH
`define GLOBALS_SVH

`define WORD_SIZE 32
`define BIT_COUNT 32
`define MEMORY_WIDTH 32

`endif // GLOBALS_SVH